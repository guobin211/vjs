module vjs
