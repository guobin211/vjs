module vjs

pub fn self_log(msg string) {
    println(msg)
}
