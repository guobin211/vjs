module v_js
