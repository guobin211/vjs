module v_js

pub fn handle_cli_error() {
    help()
}
