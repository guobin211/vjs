module v_js

pub fn help() {
    println('
vjs runtime
run js file `v index.js` as `node index.js`
')
}
